module deco #(parameter N=6)
(
  input logic [N-1:0] number, 
  output logic [13:0] result
);

  always_comb
    begin
	   case (number)
		  0 : result=14'b10000001111111;
		  
		  1 : result=14'b11110011111111;
		  
		  2 : result=14'b01001001111111;
		  
		  3 : result=14'b01100001111111;
		  
		  4 : result=14'b00110011111111;
		  
		  5 : result=14'b00100101111111;
		  
		  6 : result=14'b00000101111111;
		  
		  7 : result=14'b11110001111111;
		  
		  8 : result=14'b00000001111111;
		  
		  9 : result=14'b00110001111111;
		  
		  10 : result=14'b10000001111001;
		  
		  11 : result=14'b11110011111001;
		  
		  12 : result=14'b01001001111001;
		  
		  13 : result=14'b01100001111001;
		  
		  14 : result=14'b00110011111001;
		  
		  15 : result=14'b00100101111001;
		  
		  16 : result=14'b00000101111001;
		  
		  17 : result=14'b11110001111001;
		  
		  18 : result=14'b00000001111001;
		  
		  19 : result=14'b00110001111001;
		  
		  20 : result=14'b10000000100100;
		  
		  21 : result=14'b11110010100100;
		  
		  22 : result=14'b01001000100100;
		  
		  23 : result=14'b01100000100100;
		  
		  24 : result=14'b00110010100100;
		  
		  25 : result=14'b00100100100100;
		  
		  26 : result=14'b00000100100100;
		  
		  27 : result=14'b11110000100100;
		  
		  28 : result=14'b00000000100100;
		  
		  29 : result=14'b00110000100100;
		  
		  30 : result=14'b10000000110000;
		  
		  31 : result=14'b11110010110000;
		  
		  32 : result=14'b01001000110000;
		  
		  33 : result=14'b01100000110000;
		  
		  34 : result=14'b00110010110000;
		  
		  35 : result=14'b00100100110000;
		  
		  36 : result=14'b00000100110000;
		  
		  37 : result=14'b11110000110000;
		  
		  38 : result=14'b00000000110000;
		  
		  39 : result=14'b00110000110000;
		  
		  40 : result=14'b10000000011001;
		  
		  41 : result=14'b11110010011001;
		  
		  42 : result=14'b01001000011001;
		  
		  43 : result=14'b01100000011001;
		  
		  44 : result=14'b00110010011001;
		  
		  45 : result=14'b00100100011001;
		  
		  46 : result=14'b00000100011001;
		  
		  47 : result=14'b11110000011001;
		  
		  48 : result=14'b00000000011001;
		  
		  49 : result=14'b00110000011001;
		  
		  50 : result=14'b10000000010010;
		  
		  51 : result=14'b11110010010010;
		  
		  52 : result=14'b01001000010010;
		  
		  53 : result=14'b01100000010010;
		  
		  54 : result=14'b00110010010010;
		  
		  55 : result=14'b00100100010010;
		  
		  56 : result=14'b00000100010010;
		  
		  57 : result=14'b11110000010010;
		  
		  58 : result=14'b00000000010010;
		  
		  59 : result=14'b00110000010010;
		  
		  60 : result=14'b10000000000010;
		  
		  61 : result=14'b11110010000010;
		  
		  62 : result=14'b01001000000010;
		  
		  63 : result=14'b01100000000010;
		  
		  default : result=14'b11111111111111; 
       endcase
	  end
endmodule 